module io_multiplexing
