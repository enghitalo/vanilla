module main

import strings
import http_server

const http_ok_response = 'HTTP/1.1 200 OK\r\nContent-Type: application/json\r\nContent-Length: 0\r\nConnection: close\r\n\r\n'.bytes()

const http_created_response = 'HTTP/1.1 201 Created\r\nContent-Type: application/json\r\nContent-Length: 0\r\nConnection: close\r\n\r\n'.bytes()

const tiny_internal_server_error_response = 'HTTP/1.1 500 Internal Server Error\r\nContent-Length: 0\r\nConnection: close\r\n\r\n'.bytes()

fn home_controller(params []string) ![]u8 {
	return http_ok_response
}

fn get_users_controller(params []string, mut pool ConnectionPool) ![]u8 {
	mut db := pool.acquire() or { return tiny_internal_server_error_response }
	defer { pool.release(db) }
	rows := db.exec('SELECT * FROM users') or { return tiny_internal_server_error_response }

	mut response_body := strings.new_builder(200)
	for row in rows {
		response_body.write_string(row.str())
		response_body.write_string('\n')
	}

	// response_body_str := response_body.str()
	defer {
		unsafe {
			response_body.free()
			params.free()
		}
	}

	mut sb := strings.new_builder(200)
	sb.write_string('HTTP/1.1 200 OK\r\nContent-Type: text/plain\r\nContent-Length: ')
	sb.write_string(response_body.len.str())
	sb.write_string('\r\nConnection: close\r\n\r\n')
	sb.write(response_body)!

	return sb
}

@[direct_array_access; manualfree]
fn get_user_controller(params []string, mut pool ConnectionPool) ![]u8 {
	if params.len == 0 {
		return http_server.tiny_bad_request_response
	}
	id := params[0]
	mut db := pool.acquire() or { return tiny_internal_server_error_response }
	defer { pool.release(db) }
	result := db.exec('SELECT * FROM users WHERE id = ${id}') or {
		return tiny_internal_server_error_response
	}
	response_body := result.map(it.str()).join('\n')

	mut sb := strings.new_builder(200)
	sb.write_string('HTTP/1.1 200 OK\r\nContent-Type: text/plain\r\nContent-Length: ')
	sb.write_string(response_body.len.str())
	sb.write_string('\r\nConnection: close\r\n\r\n')
	sb.write_string(response_body)

	defer {
		unsafe {
			response_body.free()
			params.free()
		}
	}
	return sb
}

fn create_user_controller(params []string, mut pool ConnectionPool) ![]u8 {
	dump('create_user_controller')
	mut db := pool.acquire() or { return tiny_internal_server_error_response }
	defer { pool.release(db) }
	db.exec("INSERT INTO users (name) VALUES ('new_user')") or {
		return tiny_internal_server_error_response
	}
	return http_created_response
}
