module structs

import veb

pub struct Context {
	veb.Context
}
