module iocp
